// GEMM Engine with Tiling Support
// Wraps systolic array with control logic for arbitrary matrix sizes

`timescale 1ns/1ps

module gemm_engine #(
    parameter DATA_WIDTH = 8,
    parameter ACC_WIDTH = 32,
    parameter ARRAY_SIZE = 16,
    parameter SRAM_ADDR_WIDTH = 16
)(
    input  logic                      clk,
    input  logic                      rst_n,
    
    // Control interface
    input  logic                      start,
    output logic                      busy,
    output logic                      done,
    
    // Configuration registers (loaded before start)
    input  logic [SRAM_ADDR_WIDTH-1:0] src_a_addr,   // Activation matrix address in SRAM
    input  logic [SRAM_ADDR_WIDTH-1:0] src_b_addr,   // Weight matrix address in SRAM
    input  logic [SRAM_ADDR_WIDTH-1:0] dst_addr,     // Output address in SRAM
    input  logic [15:0]               dim_m,         // Rows of A and C
    input  logic [15:0]               dim_k,         // Cols of A, rows of B
    input  logic [15:0]               dim_n,         // Cols of B and C
    input  logic                      transpose_b,   // Transpose B matrix
    input  logic                      accumulate,    // Accumulate with existing output
    input  logic [7:0]                scale,         // Requantization scale
    input  logic [7:0]                shift,         // Requantization shift
    input  logic                      requant_en,    // Enable requantization
    
    // SRAM interface (read)
    output logic [SRAM_ADDR_WIDTH-1:0] sram_rd_addr,
    input  logic [DATA_WIDTH-1:0]      sram_rd_data,
    output logic                       sram_rd_en,
    
    // SRAM interface (write)
    output logic [SRAM_ADDR_WIDTH-1:0] sram_wr_addr,
    output logic [DATA_WIDTH-1:0]      sram_wr_data,
    output logic                       sram_wr_en,
    
    // Direct systolic array interface (for testing/debug)
    output logic                       array_load_weights,
    output logic [$clog2(ARRAY_SIZE)-1:0] array_weight_row,
    output logic [DATA_WIDTH-1:0]      array_weight_in [0:ARRAY_SIZE-1]
);

    // State machine
    typedef enum logic [3:0] {
        IDLE,
        LOAD_WEIGHT_TILE,
        LOAD_ACT_TILE,
        COMPUTE_TILE,
        STORE_RESULT,
        NEXT_TILE,
        REQUANTIZE,
        DONE_STATE
    } state_t;
    
    state_t state, next_state;
    
    // Tile counters
    localparam int TILE_COUNT_W = $clog2(65536/ARRAY_SIZE) + 1;
    localparam int TILE_SIZE_W  = $clog2(ARRAY_SIZE) + 1;

    logic [TILE_COUNT_W-1:0] tile_m, tile_n, tile_k;
    logic [TILE_COUNT_W-1:0] tiles_m, tiles_n, tiles_k;
    
    // Current tile addresses
    logic [SRAM_ADDR_WIDTH-1:0] tile_a_addr;
    logic [SRAM_ADDR_WIDTH-1:0] tile_b_addr;
    logic [SRAM_ADDR_WIDTH-1:0] tile_c_addr;
    
    // Tile size (may be smaller at edges)
    logic [TILE_SIZE_W-1:0] tile_size_m, tile_size_n, tile_size_k;

    // Explicitly sized intermediates for width-safe tile math
    logic [16:0] dim_m_ext, dim_n_ext, dim_k_ext;
    logic [16:0] array_size_ext;
    logic [15:0] compute_limit;
    
    // Systolic array interface
    logic                      array_start;
    logic                      array_clear;
    logic                      array_act_valid;
    logic [DATA_WIDTH-1:0]     array_act_in [0:ARRAY_SIZE-1];
    logic [ACC_WIDTH-1:0]      array_partial_in [0:ARRAY_SIZE-1];
    logic [ACC_WIDTH-1:0]      array_result [0:ARRAY_SIZE-1];
    logic                      array_result_valid;
    logic                      array_busy;
    
    // Accumulation buffer for partial sums across K tiles
    logic [ACC_WIDTH-1:0] accum_buffer [0:ARRAY_SIZE-1][0:ARRAY_SIZE-1];
    logic accum_buffer_valid [0:ARRAY_SIZE-1][0:ARRAY_SIZE-1];
    
    // Requantization
    logic [DATA_WIDTH-1:0] requant_result [0:ARRAY_SIZE-1];
    
    // Cycle counter for array timing
    logic [15:0] compute_cycles;
    
    // State machine sequential logic
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= IDLE;
            tile_m <= '0;
            tile_n <= '0;
            tile_k <= '0;
            compute_cycles <= '0;
        end else begin
            state <= next_state;
            
            case (state)
                COMPUTE_TILE: begin
                    compute_cycles <= compute_cycles + 1;
                end
                
                NEXT_TILE: begin
                    compute_cycles <= '0;
                    // Advance tile counters
                    if (tile_k < (tiles_k - TILE_COUNT_W'(1))) begin
                        tile_k <= tile_k + 1;
                    end else begin
                        tile_k <= '0;
                        if (tile_n < (tiles_n - TILE_COUNT_W'(1))) begin
                            tile_n <= tile_n + 1;
                        end else begin
                            tile_n <= '0;
                            if (tile_m < (tiles_m - TILE_COUNT_W'(1))) begin
                                tile_m <= tile_m + 1;
                            end
                        end
                    end
                end
                
                default: compute_cycles <= '0;
            endcase
        end
    end
    
    // Calculate number of tiles needed
    assign dim_m_ext = {1'b0, dim_m};
    assign dim_n_ext = {1'b0, dim_n};
    assign dim_k_ext = {1'b0, dim_k};
    assign array_size_ext = 17'(ARRAY_SIZE);

    assign tiles_m = TILE_COUNT_W'((dim_m_ext + array_size_ext - 17'd1) / array_size_ext);
    assign tiles_n = TILE_COUNT_W'((dim_n_ext + array_size_ext - 17'd1) / array_size_ext);
    assign tiles_k = TILE_COUNT_W'((dim_k_ext + array_size_ext - 17'd1) / array_size_ext);
    
    // Current tile sizes (handle edge cases)
    assign tile_size_m = (tile_m == (tiles_m - TILE_COUNT_W'(1)) && dim_m % ARRAY_SIZE != 0) ? 
                         TILE_SIZE_W'(dim_m % ARRAY_SIZE) : TILE_SIZE_W'(ARRAY_SIZE);
    assign tile_size_n = (tile_n == (tiles_n - TILE_COUNT_W'(1)) && dim_n % ARRAY_SIZE != 0) ? 
                         TILE_SIZE_W'(dim_n % ARRAY_SIZE) : TILE_SIZE_W'(ARRAY_SIZE);
    assign tile_size_k = (tile_k == (tiles_k - TILE_COUNT_W'(1)) && dim_k % ARRAY_SIZE != 0) ? 
                         TILE_SIZE_W'(dim_k % ARRAY_SIZE) : TILE_SIZE_W'(ARRAY_SIZE);

    assign compute_limit = 16'(tile_size_m) + 16'(tile_size_k) + 16'(tile_size_n) + 16'd4;
    
    // State machine combinational logic
    always_comb begin
        next_state = state;
        
        case (state)
            IDLE: begin
                if (start) next_state = LOAD_WEIGHT_TILE;
            end
            
            LOAD_WEIGHT_TILE: begin
                // Load weights for current tile
                // Takes tile_size_k cycles
                next_state = LOAD_ACT_TILE;
            end
            
            LOAD_ACT_TILE: begin
                next_state = COMPUTE_TILE;
            end
            
            COMPUTE_TILE: begin
                // Computation takes tile_size_m + tile_size_k + tile_size_n cycles
                if (compute_cycles >= compute_limit) begin
                    if (tile_k < (tiles_k - TILE_COUNT_W'(1))) begin
                        // More K tiles to accumulate
                        next_state = NEXT_TILE;
                    end else begin
                        // Done with accumulation, store result
                        next_state = STORE_RESULT;
                    end
                end
            end
            
            STORE_RESULT: begin
                // Store one row per cycle
                // Takes tile_size_m cycles
                next_state = NEXT_TILE;
            end
            
            NEXT_TILE: begin
                if (tile_m == (tiles_m - TILE_COUNT_W'(1)) &&
                    tile_n == (tiles_n - TILE_COUNT_W'(1)) &&
                    tile_k == (tiles_k - TILE_COUNT_W'(1))) begin
                    next_state = DONE_STATE;
                end else begin
                    next_state = LOAD_WEIGHT_TILE;
                end
            end
            
            DONE_STATE: begin
                next_state = IDLE;
            end
            
            default: next_state = IDLE;
        endcase
    end
    
    // Status outputs
    assign busy = (state != IDLE);
    assign done = (state == DONE_STATE);
    
    // Systolic array instantiation
    systolic_array #(
        .DATA_WIDTH(DATA_WIDTH),
        .ACC_WIDTH(ACC_WIDTH),
        .ARRAY_SIZE(ARRAY_SIZE)
    ) array (
        .clk(clk),
        .rst_n(rst_n),
        .load_weights(array_load_weights),
        .start_compute(array_start),
        .clear_acc(array_clear),
        .weight_in(array_weight_in),
        .weight_row(array_weight_row),
        .activation_in(array_act_in),
        .activation_valid(array_act_valid),
        .partial_sum_in(array_partial_in),
        .result_out(array_result),
        .result_valid(array_result_valid),
        .busy(array_busy)
    );
    
    // TODO: Implement full tiling logic, SRAM interface, requantization
    // This is a structural placeholder
    
    assign sram_rd_addr = '0;
    assign sram_rd_en = 1'b0;
    assign sram_wr_addr = '0;
    assign sram_wr_data = '0;
    assign sram_wr_en = 1'b0;
    
    assign array_load_weights = 1'b0;
    assign array_weight_row = '0;
    for (genvar i = 0; i < ARRAY_SIZE; i++) begin : gen_array_weight_zero
        assign array_weight_in[i] = '0;
    end
    assign array_start = 1'b0;
    assign array_clear = 1'b0;
    assign array_act_valid = 1'b0;
    for (genvar i = 0; i < ARRAY_SIZE; i++) begin : gen_array_input_zero
        assign array_act_in[i] = '0;
        assign array_partial_in[i] = '0;
    end

endmodule
